
module tutorial01 (
	clk_clk,
	reset_reset_n,
	led_out_led_out);	

	input		clk_clk;
	input		reset_reset_n;
	output		led_out_led_out;
endmodule
