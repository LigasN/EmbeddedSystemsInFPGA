
module tutorial01 (
	clk_clk,
	led_export,
	reset_reset_n,
	sw_export);	

	input		clk_clk;
	output	[3:0]	led_export;
	input		reset_reset_n;
	input	[2:0]	sw_export;
endmodule
