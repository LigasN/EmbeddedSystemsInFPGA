
module tutorial01 (
	clk_clk,
	reset_reset_n,
	pwm_pwm);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	pwm_pwm;
endmodule
