
module tutorial01 (
	clk_clk,
	hdmi_hdmi_tmds,
	hdmi_hdmi_tmds_clk,
	reset_reset_n);	

	input		clk_clk;
	output	[2:0]	hdmi_hdmi_tmds;
	output		hdmi_hdmi_tmds_clk;
	input		reset_reset_n;
endmodule
