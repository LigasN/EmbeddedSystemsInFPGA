
module tutorial01 (
	clk_clk,
	pwm_pwm,
	reset_reset_n);	

	input		clk_clk;
	output	[3:0]	pwm_pwm;
	input		reset_reset_n;
endmodule
